module module_top (
    ports
);
    
endmodule